`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/24/2018 05:19:51 PM
// Design Name: 
// Module Name: registersim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module registersim;
    logic D;
    logic clk;
    logic enable;
    logic reset;
    logic Q;
    
    register register_sim(.*);
    initial
    begin
    D= 
endmodule
